netcdf frc_bulk {

dimensions:
	xi_rho = 146 ;
	eta_rho = 82 ;
	time = UNLIMITED ; // (0 currently)

variables:
	double time(time) ;
		time:long_name = "atmospheric forcing time" ;
        time:units = "days since 01-Jan-2006" ;
		time:field = "time, scalar, series" ;
		time:end_date = "08-Jun-2006 00:00:00" ;
	double Uwind(time, eta_rho, xi_rho) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
        Uwind:wrf_unit = "m s-1" ;
        Uwind:wrf_desc = "U at 10 M" ;
        Uwind:field = "Uwind scalar, series" ;
		Uwind:time = "time" ;

// global attributes:
		:type = "ROMS forcing file" ;
        :title = "Hudson River of New Jersey, Atmospheric Fields" ;
        :source = "copy from latte example input data" ;

}
