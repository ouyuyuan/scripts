netcdf frc_tides_lattec {
dimensions:
	eta_rho = 82 ;
	xi_rho = 146 ;
	tide_period = UNLIMITED ; // (7 currently)
variables:
	double tide_period(tide_period) ;
		tide_period:long_name = "tide angular period" ;
		tide_period:units = "hours" ;
		tide_period:field = "tide_period, scalar, series" ;
	double tide_Ephase(tide_period, eta_rho, xi_rho) ;
		tide_Ephase:long_name = "tidal elevation phase angle" ;
		tide_Ephase:units = "degrees, time of maximum elevation with respect to chosen time origin" ;
		tide_Ephase:field = "tide_Ephase, scalar, series" ;
	double tide_Eamp(tide_period, eta_rho, xi_rho) ;
		tide_Eamp:long_name = "tidal elevation amplitude" ;
		tide_Eamp:units = "meter" ;
		tide_Eamp:field = "tide_Eamp, scalar, series" ;
	double tide_Cphase(tide_period, eta_rho, xi_rho) ;
		tide_Cphase:long_name = "tidal current phase angle" ;
		tide_Cphase:units = "degrees, time of maximum velocity with respect to  chosen time origin" ;
		tide_Cphase:field = "tide_Cphase, scalar, series" ;
	double tide_Cangle(tide_period, eta_rho, xi_rho) ;
		tide_Cangle:long_name = "tidal current inclination angle" ;
		tide_Cangle:units = "degrees between semi-major axis and East" ;
		tide_Cangle:field = "tide_Cangle, scalar, series" ;
	double tide_Cmin(tide_period, eta_rho, xi_rho) ;
		tide_Cmin:long_name = "minimum tidal current, ellipse semi-minor axis" ;
		tide_Cmin:units = "meter second-1" ;
		tide_Cmin:field = "tide_Cmin, scalar, series" ;
	double tide_Cmax(tide_period, eta_rho, xi_rho) ;
		tide_Cmax:long_name = "maximum tidal current, ellipse semi-major axis" ;
		tide_Cmax:units = "meter second-1" ;
		tide_Cmax:field = "tide_Cmax, scalar, series" ;

// global attributes:
		:type = "ROMS Forcing file" ;
		:title = "Tidal Forcing for LaTTE coarse grid domain" ;
		:grd_file = "/home/zhang/roms/latteda/grid/roms_latte_grid_4.nc" ;
		:details = "Tidal information processed from the ADCIRC database adcirc_ec2001v2e_fix.mat" ;
		:Component_0 = "K1  " ;
		:Component_1 = "O1  " ;
		:Component_2 = "Q1  " ;
		:Component_3 = "M2  " ;
		:Component_4 = "S2  " ;
		:Component_5 = "N2  " ;
		:Component_6 = "K2  " ;
		:tides_start_date = "Tides start time is 2006-01-01 00:00:00" ;
		:history = "Generated by /home/zhang/roms/latte06/tides/warner_adcirc_tides.m from data file /home/zhang/roms/latte06/tides/adcirc_ec2001v2e_fix.mat" ;
data:

 tide_period = 23.9344696552669, 25.8193416650329, 26.8683566723188, 
    12.4206012212082, 12.0000000027112, 12.658348243603, 11.9672347882466 ;
}
