netcdf frc_bulk {

dimensions:
	xi_rho = 146 ;
	eta_rho = 82 ;
	time = UNLIMITED ; // (0 currently)

variables:
	double time(time) ;
		time:long_name = "atmospheric forcing time" ;
        time:units = "days since 2006-01-01 00:00:00" ;
		time:field = "time, scalar, series" ;
        time:calendar = "gregorian" ;
		time:begin_date = "2006-01-01 00:00:00" ;
		time:end_date = "2006-06-08 23:00:00" ;
	double Tair(time, eta_rho, xi_rho) ;
		Tair:long_name = "Surface air temperature" ;
		Tair:units = "Celcius" ;
		Tair:wrf_unit = "K" ;
		Tair:wrf_desc = "TEMP at 2 M" ;
		Tair:field = "Tair scalar, series" ;
		Tair:time = "time" ;

// global attributes:
		:type = "ROMS forcing file" ;
        :title = "Hudson River of New Jersey, Atmospheric Fields" ;
        :source = "NCEP_CFSR dataset" ;

}
