netcdf frc_bulk {

dimensions:
	xi_rho = 186 ;
	eta_rho = 286 ;
	time = UNLIMITED ; // (0 currently)

variables:
	double time(time) ;
		time:long_name = "atmospheric forcing time" ;
        time:units = "days since 2006-01-01 00:00:00" ;
		time:field = "time, scalar, series" ;
        time:calendar = "gregorian" ;
		time:begin_date = "2006-01-01 00:00:00" ;
		time:end_date = "2006-06-08 23:00:00" ;
	double lwrad(time, eta_rho, xi_rho) ;
		lwrad:long_name = "Net long wave flux" ;
		lwrad:units = "watts meters-2" ;
		lwrad:positive_value = "downward flux, heating" ;
		lwrad:negative_value = "upward flux, cooling" ;
		lwrad:field = "lwrad scalar, series" ;
		lwrad:time = "time" ;

// global attributes:
		:type = "ROMS forcing file" ;
        :title = "South China sea, Atmospheric Fields" ;
        :source = "NCEP_CFSR dataset" ;

}
