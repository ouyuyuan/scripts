netcdf frc_bulk {

dimensions:
	xi_rho = 146 ;
	eta_rho = 82 ;
	time = UNLIMITED ; // (0 currently)

variables:
	double time(time) ;
		time:long_name = "atmospheric forcing time" ;
        time:units = "days since 2006-01-01 00:00:00" ;
		time:field = "time, scalar, series" ;
        time:calendar = "gregorian" ;
		time:begin_date = "2006-01-01 00:00:00" ;
		time:end_date = "2006-06-08 23:00:00" ;
	double Qair(time, eta_rho, xi_rho) ;
		Qair:long_name = "Relative humidity" ;
		Qair:units = "percentage" ;
		Qair:wrf_unit = "kg kg-1" ;
		Qair:wrf_desc = "QV at 2 M" ;
		Qair:field = "Qair scalar, series" ;
		Qair:time = "time" ;

// global attributes:
		:type = "ROMS forcing file" ;
        :title = "Hudson River of New Jersey, Atmospheric Fields" ;
        :source = "NCEP_CFSR dataset" ;

}
