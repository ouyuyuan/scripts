netcdf frc_bulk {

dimensions:
	xi_rho = 146 ;
	eta_rho = 82 ;
	time = UNLIMITED ; // (0 currently)

variables:
	double time(time) ;
		time:long_name = "atmospheric forcing time" ;
        time:units = "days since 01-Jan-2006" ;
		time:field = "time, scalar, series" ;
		time:end_date = "08-Jun-2006 00:00:00" ;
	double Vwind(time, eta_rho, xi_rho) ;
		Vwind:long_name = "Surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:wrf_unit = "m s-1" ;
		Vwind:wrf_desc = "V at 10 M" ;
		Vwind:field = "Vwind scalar, series" ;
		Vwind:time = "time" ;

// global attributes:
		:type = "ROMS forcing file" ;
        :title = "Hudson River of New Jersey, Atmospheric Fields" ;
        :source = "copy from latte example input data" ;

}
