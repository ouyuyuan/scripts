netcdf frc_uvstress {

dimensions:
	xi_u = 145 ;
	xi_v = 146 ;
	eta_u = 82 ;
	eta_v = 81 ;
	time = UNLIMITED ; // (0 currently)

variables:
	double time(time) ;
		time:long_name = "atmospheric forcing time" ;
        time:units = "days since 2006-01-01 00:00:00" ;
		time:field = "time, scalar, series" ;
        time:calendar = "gregorian" ;
		time:begin_date = "2006-01-01 00:00:00" ;
		time:end_date = "2006-06-08 23:00:00" ;
	short sustr(time, eta_u, xi_u) ;
		sustr:long_name = "surface u-momentum stress" ;
		sustr:units = "Newton meter-2" ;
		sustr:time = "time" ;
		sustr:scale_factor = 0.0005 ;
	short svstr(time, eta_v, xi_v) ;
		svstr:long_name = "surface v-momentum stress" ;
		svstr:units = "Newton meter-2 * 1000" ;
		svstr:time = "time" ;
		svstr:scale_factor = 0.0005 ;

// global attributes:
		:type = "ROMS FORCING file" ;
        :title = "Hudson River of New Jersey, Atmospheric Fields" ;
        :source = "NCEP_CFSR dataset" ;
}
