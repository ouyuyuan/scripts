netcdf tides_yellow_sea {

dimensions:
	namelen = 4 ;
	tide_period = 8 ;
	xi_rho = 82 ;
	eta_rho = 82 ;

variables:
	double tide_period(tide_period) ;
		tide_period:field = "tide_period, scalar" ;
		tide_period:long_name = "tide angular period" ;
		tide_period:units = "hours" ;
	double tide_Ephase(tide_period, eta_rho, xi_rho) ;
		tide_Ephase:field = "tide_Ephase, scalar" ;
		tide_Ephase:long_name = "tidal elevation phase angle" ;
		tide_Ephase:units = "degrees, time of maximum elevation with respect chosen time origin" ;
	double tide_Eamp(tide_period, eta_rho, xi_rho) ;
		tide_Eamp:field = "tide_Eamp, scalar" ;
		tide_Eamp:long_name = "tidal elevation amplitude" ;
		tide_Eamp:units = "meter" ;
	double tide_Cmax(tide_period, eta_rho, xi_rho) ;
		tide_Cmax:field = "tide_Cmax, scalar" ;
		tide_Cmax:long_name = "maximum tidal current, ellipse semi-major axis" ;
		tide_Cmax:units = "meter second-1" ;
	double tide_Cmin(tide_period, eta_rho, xi_rho) ;
		tide_Cmin:field = "tide_Cmin, scalar" ;
		tide_Cmin:long_name = "minimum tidal current, ellipse semi-minor axis" ;
		tide_Cmin:units = "meter second-1" ;
	double tide_Cangle(tide_period, eta_rho, xi_rho) ;
		tide_Cangle:field = "tide_Cangle, scalar" ;
		tide_Cangle:long_name = "tidal current inclination angle" ;
		tide_Cangle:units = "degrees between semi-major axis and East" ;
	double tide_Cphase(tide_period, eta_rho, xi_rho) ;
		tide_Cphase:field = "tide_Cphase, scalar" ;
		tide_Cphase:long_name = "tidal current phase angle" ;
		tide_Cphase:units = "degrees, time of maximum velocity" ;
	char tide_name(tide_period, namelen) ;

// global attributes:
        :title = "Yellow Sea, Tides forcing Fields" ;
		:type = "ROMS FORCING file" ;
        :source = "OTPS dataset" ;
data:

 tide_period = 26.8683567047119, 25.8193397521973, 24.0658893585205, 
    23.9344692230225, 12.6583499908447, 12.420599937439, 12, 11.9672346115112 ;
}
