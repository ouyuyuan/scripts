netcdf frc_bulk {

dimensions:
	xi_rho = 146 ;
	eta_rho = 82 ;
	time = UNLIMITED ; // (0 currently)

variables:
	double time(time) ;
		time:long_name = "atmospheric forcing time" ;
        time:units = "days since 2006-01-01 00:00:00" ;
		time:field = "time, scalar, series" ;
        time:calendar = "gregorian" ;
		time:begin_date = "2006-01-01 00:00:00" ;
		time:end_date = "2006-06-08 23:00:00" ;
	double Swrf(time, eta_rho, xi_rho) ;
		Swrf:long_name = "Short wave flux net" ;
		Swrf:units = "watts meters-2" ;
		Swrf:positive_value = "downward flux, heating" ;
		Swrf:negative_value = "upward flux, cooling" ;
		Swrf:wrf_unit = "W m-2" ;
		Swrf:wrf_desc = "DOWNWARD SHORT WAVE FLUX AT GROUND SURFACE" ;
		Swrf:field = "Swrf scalar, series" ;
		Swrf:time = "time" ;

// global attributes:
		:type = "ROMS forcing file" ;
        :title = "Hudson River of New Jersey, Atmospheric Fields" ;
        :source = "NCEP_CFSR dataset" ;

}
